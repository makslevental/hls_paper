always @ (posedge ap_clk) begin
  if ((1'b1 == ap_CS_fsm_state209)) begin
    reg_1608 <= fu_1076_p2;
    reg_1613 <= fu_1082_p2;
    reg_1618 <= fu_646_p2;
  end
end