always @ (posedge ap_clk) begin
  if ((1'b1 == ap_CS_fsm_state209)) begin
    notlhs17_reg_1608 <= notlhs17_fu_1076_p2;
    notrhs18_reg_1613 <= notrhs18_fu_1082_p2;
    tmp_8_reg_1618 <= grp_fu_646_p2;
  end
end
